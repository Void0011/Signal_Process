`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8HN++j8TCvG1mG+mn/45Jt0YB0PFV2E+H5+JLABBfWOkY5e22U41RTX7qT9fskKG
aW0Omz7sz6UpESXk9wvuRrDw/WseXDJHmf59DDKiu/6oaErZgdECHAQGY719fgJz
iS1c1QDL+5FRBQJq4nwx4t1uvfl2VrtZ0BzK0NrlpiI/vXliInIpvoIb0jwoepsQ
jL5aDh6snfr78W581nWNwNRRFPU4iTUhsRC5oLgshf4h5HA27phXsGKX1YaMWNRh
cy1IND7xEX4BpHvIgxnMsQGhWfk6S4biEvDjAREpgsX013ke+4bufvXTx73qUbwS
rmIj82sF6EW7Pk/gS4B/fEu0EfwmYkqaQQkCTJBqPBoVH0MzqSQru1h1375ZYGJ/
4QRiIdCwLQA+u9Xtv9vf2V//d7Xz6CzCszdrZlLNvt0hjcKKq3nocUE35sVLJx2S
DFb3JFA5oAoF6LWeYoYfzroiMnbs8DD865vaqIjwyK+u69mg/cRPV8OWc6T2ALYL
qHqm7JRCB03fRtsiIJnSYUUWglClhbSlf0qAY8L4+EAitxJrkSsPygGVLCggcpQg
G32jCBzu2JlRbJTLy4isNtoWv6vmHNeTikKLwWVdmfn0SsWbvNF4uZ5ei1NTMYRl
XVBDavommEuyaoqpn0RNB1957p23B0MTquIpu0nRppU+stOKY9NbvQ2PHE8G8n9h
ue1bSZU8/8vwwrxszaKGHKBpNoj+Wooi/oOzYzwp9p+ZaSLJ9d8U2cnJ5qSKSnC1
52ZUKNjBpp+4wEU4327FqxP+mWgLpQyTFa06cs/hG1UzABZMQdI4hf61D1OgJ7rQ
G5AnyjCIvQkb05rIx0FmdkHQS7048a/wLoJrUBMKUg2IAZmKaWEa+noUlJ+eKKD/
OjIyzPJ29MFHwyE5kNqbdEz0nxZpPN4ej7fdZ9+pDs18hVtFQvS/egKVjNlg1050
KaZvRaXg/rB3A+5faBiQ0TLqEkjiU7/iFQceNfkD3ApjTq66CvplsyOjX6vFn8pI
PB0NNKcDoH+Q8nKIPBhteiCow/yh43X6CqmWztx4/uKT1Tg/qzENgeTykaMdTR5Y
`protect END_PROTECTED
