`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kJu+tXHdScG3CxdoGoyZChtADzndG4ZNy2RqKpH4MoLGeM8awHpda4RggriDPb/c
Zb7JOKAGfSjZ4RrlWnYV+9YWO6h5LB1Vs6k9Ef6ewsgQ56bLCwZ1nz6hRo4OxW5K
Axgbi1KxOHUJj0oIG21NyL574OGUxXULEivKAt7fttnisl7Sxhb2sp8wsz6Cg3t6
IJmDhpjY887Wdz6xKSD0LTT7LvZD/rTb/7183p13VHkF/6FC9Y7JLcwg094ZVVCJ
4Pq7jHhehCvfIWc1FfHiTh2MDl31HwMy007BhnPL0stSiFv9HpxCF5U2cXXjbzO/
jyBy7I2UufOhRr672TRA1dZxBOWrd2rk5Rh3lDMrGUpnwJDji7jUuCHbldQaufy1
XF9E6bULa9tXKQhrNwmvcKu1JYateorAoutYQ4MEgzN9j6C7MafSVBOGYgmlYT3v
Ljdxdk38jB+Isk1WgPevfF2acKaNgdaEcztBosdGyospyC2fJNCM0O3rM83gEd0h
S2PN2M/IhdEXIwb/cJgeJtszxkfcuTNJsbBFgf7/0q5LVkGWpdC6ZHvW/+dt+pGq
Cwic8hbI97IhDc2nf2FHb5O3KDORCkHuzBP/mG+gMvkl9xvvRE8MDBw5+yzUvE44
aHKGFXJ/lQocmSGOdsR0zpMfakUvaL35FPKjmWX5roWwBskrc8cq7SHBckFsA4tC
497r1jHOmxc6j5KfK5p7+hSAvZzgNURJpYTbuau778DWeP6JqERtwKCr9SCyY3Ik
RBbuqelVdqw3U3oIZfgB+5M4Rum10dU1aB3qdIZ0W2i3ycrXJRJsI4yMhNFPVkgd
BCKkGT4FJA2nYGt863vqfp0ZSd4iGd/KELN22/kMyBWnCOXSc4IMI3Sc3UcjwCIv
RJ3iIOaMfiZVEmC+nlEumg1jfD492CnFjFUk5wuGPcO/gMzKNhA8dOZYQOoe3Nh4
XtKXOhj6dTXyRGFdVlFYTnzVUWtPRmbUzR/oBjiTuqQH7rvcn2vdFwzAH++BY1Lu
LFfs8kxzRtijfdyT77m2xoxnu1+sSjkk0Pfv63YGJQxY9BMLXqvSJIFglXC7S6Wt
hYyhi2X256mRuFpFfDsRZr8WyvG21GLghxFncYPBL22oj5qsDSo8fpUO0Hd3EnP6
b+eSOrGDQ68PtDeCa5p5f8sRdGulqp7lzNoIirhbR4NnZtsq/+htUumzl3Q4CxrO
FFtX25RswNLRw52LFdpNh+clHNvTKKD5YuTC/EtRHqpZaeQy1oYzqzLqf6sVrlkr
WGw5tLqnhgk9bIySL8DCMFYKvbikcqtNUZbnf2UT2M+C0icznaXR55G9TuRlIM0a
KR/c7NsDwCX0Pe40TmWCYYMiBD/3xkfTr+nsIXlsqQiSjJC3J/a5kYJpLtpZggXp
6ZDRUHdiyryFKr1Nbcku3N+Ue2T3+tHlQasPu1brm2HBphkXLjqm5l1ooHJ9WKLx
peqGl0N8F4tQUBTzFBBygSKe9roIzA20RQZDw9+akWsrvXIz3KC1JC+HdpI2U2tH
0FD0eqWlY3HQPwIBqDflY6vx2JahSAxjhnKLNlz+/e53mXhUTJdR4i5/7sED4+fr
mrtI5RJwIRqs/lOi1Lz6IGrXzkvJZ9ERJlOuGJ5p7jBHmbfbfPQ/ik6C/yjl7W8s
Y48lI59lOnKv9VOsNTQljWikt3FGReKQqsgm8ssGNEGt6n8tvVp93EoOM3QJyikY
8ye6SNqqYc9D7frojjYEFoeuEDRBUHWaDkCC8yQeTQ07USBvg/so6jTqLoleyYOp
kTrMSOQmGyRIIdwTDCwFU6xRAfgm+ssUlF/L3yXNidEY6T1Za0pk1WvXjmLckpL7
mvAtTwUh6++u580wUUoY4pPiw2JtkBjbYE4u1VzuwTZ9wzzjrvKl9kU9cjYphz7a
0LOLzxchEoqGSgcKFsxkUmdf2ecNOteVMfSvJ6mkkxkwvj34+0Kj09/uXPc1p/gR
YyJEtPVtBKAoqA3QRKGzJYhpuYb8M7qjMNx5ZvNDxPplvUWGA2GKky+u/kpG07IS
`protect END_PROTECTED
