library verilog;
use verilog.vl_types.all;
entity A_RAM is
    port(
        clk             : in     vl_logic;
        rst             : in     vl_logic;
        initial_en      : in     vl_logic;
        datain_re       : in     vl_logic_vector(23 downto 0);
        datain_im       : in     vl_logic_vector(23 downto 0);
        wr_en           : in     vl_logic;
        wr_add1         : in     vl_logic_vector(2 downto 0);
        wr_add2         : in     vl_logic_vector(2 downto 0);
        datain_re1      : in     vl_logic_vector(23 downto 0);
        datain_im1      : in     vl_logic_vector(23 downto 0);
        datain_re2      : in     vl_logic_vector(23 downto 0);
        datain_im2      : in     vl_logic_vector(23 downto 0);
        rd_en           : in     vl_logic;
        rd_add1         : in     vl_logic_vector(2 downto 0);
        rd_add2         : in     vl_logic_vector(2 downto 0);
        dataout_re1     : out    vl_logic_vector(23 downto 0);
        dataout_im1     : out    vl_logic_vector(23 downto 0);
        dataout_re2     : out    vl_logic_vector(23 downto 0);
        dataout_im2     : out    vl_logic_vector(23 downto 0);
        initial_flag    : out    vl_logic;
        read_addr       : in     vl_logic_vector(2 downto 0);
        dataout_re      : out    vl_logic_vector(23 downto 0);
        dataout_im      : out    vl_logic_vector(23 downto 0)
    );
end A_RAM;
