`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WW6uOFnYr4USWu2iICyNNBVT7EbVGUsQR9imtAi/1EHqP90Xgq/dEqyfpqt1VkNW
UfrDdg8dtgLMJZ2qcIQnAYVt20oriKcDs7DEr6TeXzrItm+5tE0UbciGRFDBrGOG
v0oaGCCq+/fh2Jlnctz/KiVE7GruGxIoijr6zRA+G6Sri5EXLvqmrO0jd0W7zq/i
nlqcNUJY1TfkFBxzt4AcQPLyrkN9c2IB41dqo4wb9Wyps9FnkfKp34iludXMrbAV
LJV4Jq22Kd4RwvIaCh1qKIhj6mEr8b/gsUwqTa4f2fuG17JrpWelh/MDygPayHnE
NSwJxuBz0xv3iv/YmM1C828wlyz5sPdpQV2QIwGGNhV99hcLwKsWcAG4CSoUKqvY
gL8S+x3PkYgRZi7fX4E/CAm2gJbTkLUswAxPZoS+gui/L06IikHb3MtzJxBZ8tq9
Bp/tclqmqqLT/gRlWs3Dral+6N1CUxhenuGmY3OUEFiSeLjYX+7lygataBGq+j8k
xElzlfOpC6oDuvlUNsueSgDWXVek1sb4HimHr1NraZ5bXdO3EqUX3AlaaV4cruz4
sldjA1enXy8dpRmZLwXyFk12qO3tTIuOPJ79hWG7WoLDUdOSBiRpncv222ODMLu+
2tNqOBvrUPYbTe0iBxIqZdUAkecOKjdWIx9z2hXgn1ca06xQZFzwQx9kKbTeDeIe
85PlLrdLWRPqbBuf5KtXrH2ORR+5+OfrpUB3GdyMcqUP9L3j/fM+M6KRTMGi18k/
hXf4CKbKw2FJtH8WiNTQvsKYzx+B6hN1cxWKk3yt02E5tOxf6F/Mx9Ihx486XJUb
9rZUsdkWwON/z2KmYHAJuzTIEZ329XuoEgiT0xGPOoM7sYlADGDg3A9VZusynp3K
h3v2L/p716BuzINvZ+jbeR9sRThFw4ExziTTbzKxuAgVy9YeTnpp8eRvDgDDx4r5
17fL2o9Dyvd11MR/+zI4RxjqbR9/umCZNhBVEeON5wMl9rHOaX/vXg+6n8Rb0Rf/
9qTtwUw+1JQ/AXmV3keNXyA8oAdIm77LsPrnzR6Be3fJ4kaSfUN3RXCT3LZtdV/k
IYpgPtp+H2oX5MvQ7eTgkA==
`protect END_PROTECTED
