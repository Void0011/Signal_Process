`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L+pKfDuJdSj5X5LmOK4o1ZHpkr2u+t2FgkRspuX4H6PngzbiHk0sw2PZdrP6zerl
rFMHpT8WF8ptplKhMQRA+1pka6VDlHfeaJG2giva0aEqWF7QSaSOpX7FRHsK3REe
/nkJkIpNRinILExSe0bCZyzL1Z/7AgbZjy/BlApHWCoNFObjji1V5ZRfHB8m2Bc1
MlVmFDISYoS7kqyp81cIsAeFoUV0qt7c0DbPe8QCOCZSARVNrS+/SKTw+Npmby0a
BSOyTha16cbiJZ+GyWxt9NsiKNlbSSfHtedwJqPJCnkZdPm07Zubsz1d0BOD8cZA
2JKmdShdABc61YUnd2eg6Av7X6ITZCn0sbrzb4A4zmcTvcCVNjhcvlXjyeikV6QJ
x+uvRaxu5ZHAO+3Xc+7izSL9HdawI9SKVDTlpQQjilMFPclG44Kh8k5EfgQbynM2
S/6Aj1K/rbpVI0S2L3IDS4vuvsLDB80wPKI0TzV4vzI65NveiEyCBOJIApadySzY
IpaRUbvjAFvf4f1zF08YdgNPJgOB8KIFl+OYrUpywhzqV2UOTjjOMXZcFhSytfXd
5uVOFkTzqdpDhNNnjqS4QjSC3BYSJnhZkbpt0RtZZCo=
`protect END_PROTECTED
