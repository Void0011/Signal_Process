`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1nLycBtfD4bClHTaDeD4R/g15Z8h7yOkq6AgOEuZgU+Rkp7aqh6gA5TJCm69zbCQ
Pao39aLpa8pLPJDo0IKGqVNUDnGpS4Ak8w5YzGLh1Ajl51Bg/9+PeTdho8Vw+wVr
Y6U0l6XZiRi7qfkI2EWA3kah2nEzoH+ZY/j3dUfwCVSQQPcAfSq+NthywJTjwzok
yOvUkzI5KeACRVvFOsH7xSMunJOAqZws6uhqi820+ezeA7gOTFOr9sFFB1f45wXI
RRGLbS4YUCJx1QQTAjazSYlUCytQzYZnjLXYCWGVruQCn9z06/MdhjDniNG9azXM
xX4vOoVRb8pAV0eKhM35o/TaXhYA4QVk32/o8cYfriU/TLGgCFigU9IA0qVF5KmG
R8H1yUbGEgvujTHjF3dtCUhYc10JbDWS1sOB0gSWT4/vbKgCKyqR4p+H5e/o6as4
CHgBHQNH8uCccE3wtNlNIJLIzHSKJoBtvNFwBOtVRG4I4Op0pCzGf6jO1MxLLqgT
uO1uKk+GMMxRZ8C9v1wa24E8ngypApUG5cyjDCy6y4ROv1AQ55RE0A2NcEDymsY5
85yVjmKtydfZlEWRBP0zzfWBMwr2rJ51jiycqLoBUYCg+KtJSZIGvG/DhJzMQQp8
P/2Ogm4mHKHFy3UxTznilC6TgETQRGsq7/8BiRhCyY6BEopseNYTSmN7opKclp50
4e8PDzj9XkTM5krIp5hLXd531vWFwmz/gpttMXeYvsg9CQjxI1ZevBN0/nqYIV1I
OZYKEHsweD3utNJt3cCVl3OgfCDj4aja4P2q/OWhPP2UfqUJ/16YUpQvOO6IM1OG
K0VaonWmD6IocIQcN+8i6pt1Cof0QeFibLMMOPFJg8Q=
`protect END_PROTECTED
