`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
njaGGewvJf74bwJqkzwezaoMhnMYbuqGi9/5IY68bnqGSxCv3ROAM9pQpZJ7SurW
bN8lSnHKXm12wfVkf/vDNY2m5hjPc+T6SnIc/vL5frI74RmFURxNZE1VJ7vMXT3m
EbU8LCE4V+Mypgj+6b2l9u21gfEtsVwz8nO7/syOo8g/2KvHVfmTLX9wFrokKaQ+
NLXWp6GrZINpaKIiJnDnN5+Ijl8ZjELA/AgvgH1hsakFi1eAd1QX5VLV6Uu2srgD
ohDK8dJpWXSfiiHWl5GbDcI0KqYFRMXFNWDoQ6tPWD7CN9VoHou4WGJK+xZRpq4b
RSMdS3DMbxisP1lfV/yVUYzTaKE57CPRip5kfDZs+XysL4Svu1/HdL/b2Cdz/5Jf
MV5Lh2YDoFJDGdXnU1dDznZmebCkYAR4KuwyAF1boeIFJk3BIcbDdVeZXDLE8pOP
wpe+uNAK7XH7UCTjv4yNdtSMuZX9GIopzk2bTHbT5tRWkFZ6dqW5TwWWxM2FL5z3
9CnfXLx4Kb/Yt3jZO9LK5c+aC4mqzGO3eAzS2cIzBW7deYCU6L428xluKLfNwstG
2PaPmlVTvuI5GyMRojldfXdaH6UiVKBAxPjH4usRxutdItdEy8ysPCeEtVrbrtUE
GlwHgf175Ck6LX6MjUZSEe19nQfGMWeV70YfbDh6BDDrQLSnvkE4LmTBbIvBTduP
LurB2LSgUWBCQYmjEJ5ttwKdg8Kxm/qiGQrKsCpi3T+b6OnuIi8kyk01m3UdhrF/
P38ZO+RyffwiM9tsiuVQcN1SPKfRzLdi6k4spFNdW1JiX6HjqLzfc9RuKymdIWO0
3XwGanZUux8PTB0Fwk2yipcMjdTKiF3e4k8vMHsH5DVLeHrLHiS9iSPjDdhbryYo
Ll22W2qls6UKWlpd47xW4uIVxybnH34ErmBOZ8GBOqpao+4QuVNuXepRJEWWTR/R
PGWdmGPVGgf8ImNJSMKX6fKls83udzzEWotB1nKF5XIPv0e3rO0CAIAiszDWfqTO
CzBc3SL3/UZn0GsIPnYbCFuyqNPtrgA9Nog/fRvPcoGBs8nPRRbD1N0pCk7d4Sd2
qzAkxBqLnkj6HKE2Ab5tONdUmtebMzwN9EJAv+L7gE2zKYoauwkvIT3AW49l7xj7
WhG1ko/Uc3MTbBW6jmHCuq6euCfl5d21LgMlCL+oBQT+x1yLx14fm0MALjAyIGi5
8DOEHkkrpiLfNEQnZUyMayBWaut53wesAMiaEnllqVTF8vciDzySEI41EHRQ4+9f
yx+M/ZyvRXAP+A8VK8FXMLZonjZCUwYE4PfY3uIGQzjRDnv4ASPuab+ghgAz9qd2
`protect END_PROTECTED
