`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6GcKF+k6uhvDwmlnrP1jQ9LQN/rOGptPYXkIVVGtHD2c0fxhQ7doW8tUqAh1sOZh
pu1XVgidg4aUJnQmbp+KlQmxvqRc03QRrSy2vLU4nCl4a9KSnq3Ip2OqyWkdCq68
ER/kVR+db/n8Y0sevDsZOKdSXT05hrDpvT1qrZwmkLllGExg80qgKqZvqPyne99c
OIcXa66AoslnbSZTP3KHD/Ig9dsTLLamTyxwAyA5eybqyEE73X9ul0FkCXFSmOec
9j/Bi43t4pM4gRqCVatrToIhHsdO8ndz+NOaVQo1U0kWTVwf7rWLmjK6eiCmOIsX
0cYh1qpBjdAi1pLPFKGEXcZbr1CPY2CyIyV9NdImy03qYvJ7b3Z/drhHoUXOu6Sg
JmYCeOLmJ+cBbr6Do0SBn6QE0K5vL82a2S0iP8UszXGE4Z8xYeR/4BNlsotJUPy/
8VwnRyWIuWg/mhbYWQKieWLKIhsdZYcTGUgN/UefumgexXLLRYrICEvpDp34psud
JCz4bFcIxSUHeFAwicV+9xJr0q1RniYPRItIeJh9R0xV4gVluoyymTeO0VfiOof4
QqAE8oa9LdMLmBND6b5FSjjJ/QgrhU5K3ZUoiSP0s2yqPTDCAlcswdiJX1+sWQbu
nBCEaN8L2A6wnlNnMuMTUMxWWfcdM5IDRbNEuN5zgiurpJB0m3+6MjduWQDfW0VN
aBJrHhF9vjiyXjPUuIN2G5aeQtdzt/OKam/qtOMIekg5r+2+bTkm34zyTqdvvn83
qrI+kaTP3IoXm4OFMRiCU0bqkfAiUL57YY9y86jxnBL5X8tWBKD1PeyvyFmD/7tV
st6zuZH9mTg6kGlPjb06oEJIk4NLOERG7rG29RDQDBQ=
`protect END_PROTECTED
