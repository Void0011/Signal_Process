`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ov3fzItbvkfhQ2A5A1TtTILy5B2LkdXCLiyL9XVMxRmLmfR2IW125lzCPDGAeGvO
pTws/c78sZ7VqFcyUdYTtUtA4+UYnA5ZF0COsoRp3naB8b6hFOW0KIueFhRD9GUd
fVVaCGxEdm4kxay8F5PI2OW5adm9SExpTA/GTBme8o5O6HVWd2VYy3qTZLvfN2fF
/sZ0B+iZNPt8EUKGUuJr7BDzGD38suJCrxcnEeGBaV3FwGvk1wkZ4Y7wrdcV9fgG
QbdrA7atwMFymbB6y/NWDgjbT+1+T7FIhKZRAgZeymlX1LOTPlg/XCRD+AQYW+MK
Rn0JWDEOtYIQ9Q9p/OIuYF6tUh9J2Zp/ovU059GAo0hW9Hmw8lKCAekLNwcOncIb
Fpj3AJXLjnpaeyTni0/qYNOcYpFYFLiwJEmLMHIPYjy6Ej6+pCd1Uw31bt5Ps7ul
AIbt0ryerP0CH7725XeFfwFb1Ms2G+PWrhf1IQaYP11GczJ/JGkFucEiaXI/ENLw
Qtkhfi4duYDEfLwvP+3iAcI8tvywXwEtl98Gn0fRMoP3PgLOoX5QrId1BuZ/cz/r
vcMSxsiQ7+X9HsSiQWdcOjCSxWJvcFmDO29UiF0fz0dSvuGfvozzOOrnks7G4caT
PeY4OQpfxYtWp4eOjJcPPVeuFnppxBSdnwuZNT2klK3O/Eyn58vXbP3aiMfq+sXO
`protect END_PROTECTED
