`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hy+PqWtAO1bxIehwiSwqNvMQ3CAQy1yiY/47qYuW0JiaKfFdgcG8XNoZ5klEVM30
YO5F6q8k3edFgzFrvmarNWGDic2PS/rpTiqJkNcIpYe5eLqoZzD8F/JMpYYw27GV
3d9arNwJQOayjLV1stEpMErJ1sEpFnjqnCxFP4zifvERUq0KYQAMefJuHlAbNtwC
yFkPrOsolfI+lvW671b0WbkmOqUCuLBRKGWxGRH6kLdjTyxDspfK8PaKdSyghFI1
KmCaIP7ZWrK8ebFjxN46T8UtvyyAkgty0U/HXwCnKqijH0kI1IXnbxZFTAb6ddrf
Rahi6fb8nfx49TU+m0fO2JVmkZh0TEC5svtlTGQjZQcGyL+L2JGWccT/2NPOJoej
FlS9R3KhtATeqe3LNEpLvq0tXRVx+tIpgFA2diSnvRCru1ZtKOsXIQAp1UOctr4v
cf6EixRSJBZWwWLSmzjrXqU3pwNN1GFzli+qYtQr/4ty0rNHVIyuKqXVwojiBsO7
qXIbMDP/kMnC3ISeK4tSh6F+StgLzDK6hOYBDCE7gjk9lAmmGyEbElDsWRkAyiu3
VyRZkzfuXlLrD2+BKihkHICVZwzJ6P3qvXg9h+GRc6hoG3ZT2t1V1J9MTC9dgsYw
OIF7XByom2GIYBsZb/VDow==
`protect END_PROTECTED
