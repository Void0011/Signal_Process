`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k+qhIEzWBoB0W7SKjBPfg3S0S3vb1H3/GaVnrNoW1JJYZUW/dp1yNo5OGj14MTx7
RoUddJ0u5i7/732xJ/WSq44izuPWDW0fJHtQMwdi1jp8Mbb/MDa2GfoRlI2Edt57
CLTeSzuACuyoAmoIc0W7/CyxUcO92oQ/QT9yLgWspt4JpLjuyyzcJc1/Klq6+3GE
d9c41m3gFObkAGUSnc/MkX24v3go8FSx01fR5ty5vxohN/v1CelsrRQAa3zshU37
vy/a9Lo3whGzawkve1wNsI74BNj5GhgjpHENu9/zlqu25qPiL/Z5JzpLhN/yrmB2
3/hVS2VaTf9yyOBCxk612iXWvdr2wUcF/wy8T7bKG8uv6Bark3e99kqvZlReEM2X
hfTmwFyvY6RTwMWtqmkZXUFiG7viJiP63yIe/LQZY6BiOFOAmAS2Tr+5ZrWOptQC
2N2YbJuolZwoa6+J4xY32xWtiYCiH1uk1Vjz9p3IXzQ9ggKcuRJmjSL6qA5PmW8u
7NXjKu/xnaGZusTjDCajiY11Ye9Cc/ZfBbCa8I5rYkPJB800Bwye9YCBpUX76sqr
IpAj5xLWKDlukK55j6NBpfr8wJAiJYleg64vYR/+vPfbPcChpF7LtJcN1/aDuOPB
HQtdCKf54zQQ0Eg4ZK2HSKe1iuWEG0AOjmQlFcq2c6qYHPJVHJEbc/NXxgp36NC/
3me44c4tlpcQGBny8vvQazNlZZdQVIE+5fpx7jP1s+g=
`protect END_PROTECTED
